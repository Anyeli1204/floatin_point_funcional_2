module contador(
    input cont, clk, reset,
    input next_row,
    output reg [31:0] next 
);
endmodule